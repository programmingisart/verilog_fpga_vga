module vga(
	input clk,
	input rxpin,
	output reg r,
	output reg g,
	output reg b,
	output reg vsync,
	output reg hsync,
	output led

	);
	
	wire pll_locked;
	
	reg clk_25mhz;
	
	reg [9:0]x_pos;
	reg [8:0]y_pos;
	

	wire pll_25mhz;

	wire rx_byte_ok;

	wire [7:0]bytes;


	reg [1399:0]datar;
	reg [1399:0]datag;
	reg [1399:0]datab;

ttlrx ttl(
	.clk(clk),
	.rxpin(rxpin),
	.out_bytes(bytes),
	.out_byte_ok(rx_byte_ok)
	);

initial begin
	datar	<= 1200'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010011111110000000000000000000000000100001000001000000000000000000000000000010000100000100000000000000000000000000001111110000010000000000000000000000000000100001000001000000000000000000000000000010000100000100000000000000000000000000001000010011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
end
		
always @(posedge rx_byte_ok) begin
	datar <= datar << 8;
	datar[7:0] <= bytes;
end		

 pll pll_25 (
	.inclk0(clk),
	.c0(pll_25mhz),
	.locked(pll_locked)
	);
	
always @(posedge clk) clk_25mhz <= ~clk_25mhz;


always @(posedge pll_25mhz) begin	
		
		x_pos <= x_pos + 1'b1;
		
		if(x_pos == 800) begin
			x_pos <= 0;
			y_pos <= y_pos +1;
			if(y_pos == 526) y_pos <= 0;
		end
		
	
		hsync <= ~(x_pos > (640 + 16) && (x_pos < (640 + 16 + 96)));   //96 clocks
      vsync <= ~(y_pos > (480 + 10) && (y_pos < (480 + 10 + 2)));   //2 clocks
		
		
		if (x_pos < 640 && y_pos < 480) begin
			r <= datar[(29-(y_pos >> 4)) * 40 + (39-(x_pos >> 4))];
			g <= datar[(29-(y_pos >> 4)) * 40 + (39-(x_pos >> 4))];
			b <= datar[(29-(y_pos >> 4)) * 40 + (39-(x_pos >> 4))];
		end
		else begin
			r <= 0;
			g <= 0;
			b <= 0;
		end
		
end

assign led = pll_locked;

endmodule